LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--use ieee.fixed_pkg.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MULTIPLIER IS
	GENERIC ( N, M : INTEGER:=24);
	PORT (	A : IN SIGNED(N-1 DOWNTO 0);
				B : IN SIGNED(M-1 DOWNTO 0);
				EN, CLOCK, RESETN : IN STD_LOGIC;
				OUTPUT :	OUT STD_LOGIC_VECTOR(M+N-2 DOWNTO 0));
END MULTIPLIER;

ARCHITECTURE BEHAVIOR OF MULTIPLIER IS
	COMPONENT REGN_EN_FP IS
		GENERIC ( N : INTEGER:=24);
		PORT (	R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				ENABLE, CLOCK, RESETN : IN STD_LOGIC;
				Q :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;
	SIGNAL M1:  SIGNED(M+N-1 DOWNTO 0);
	SIGNAL M2,M3,M4:  STD_LOGIC_VECTOR(M+N-1 DOWNTO 0);
	SIGNAL EN_0,EN_1,EN_2: STD_LOGIC_VECTOR(0 DOWNTO 0);
BEGIN	
	EN_0(0)<=EN;
	-- STADIO DI INGRESSO
	REG1: REGN_EN_FP 	GENERIC MAP (N+M)
							PORT MAP(STD_LOGIC_VECTOR(M1), EN_0(0), CLOCK, RESETN, M2);
	FF1:  REGN_EN_FP 	GENERIC MAP (1)
							PORT MAP(EN_0, '1', CLOCK, RESETN, EN_1); 
	-- PRIMO LIVELLO DI PIPELINE
	REG2: REGN_EN_FP 	GENERIC MAP (N+M)
							PORT MAP(M2, EN_1(0), CLOCK, RESETN, M3);
	FF2:  REGN_EN_FP 	GENERIC MAP (1)
							PORT MAP(EN_1, '1', CLOCK, RESETN, EN_2);
	-- SECONDO LIVELLO DI PIPELINE 
	REG3: REGN_EN_FP 	GENERIC MAP (N+M)
							PORT MAP(M3, EN_2(0), CLOCK, RESETN, M4);
	OUTPUT <= M4(N+M-2 DOWNTO 0);
	M1<=A*B;
END BEHAVIOR;
