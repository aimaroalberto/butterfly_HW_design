LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INCREASER IS
GENERIC(N:INTEGER:=4);
PORT(
X : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END INCREASER;

ARCHITECTURE BEHAVIOR OF INCREASER IS
BEGIN
Y <= X + 1;
END BEHAVIOR;