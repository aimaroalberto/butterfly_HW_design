LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ROUNDER IS
	GENERIC (N_IN : INTEGER := 49;
				M_OUT: INTEGER :=24);
	PORT (	INPUT : IN STD_LOGIC_VECTOR(N_IN-1 DOWNTO 0);
				CLOCK, RESETN : IN STD_LOGIC;
				OUTPUT: OUT STD_LOGIC_VECTOR(M_OUT-1 DOWNTO 0));
END ROUNDER;

ARCHITECTURE BEHAVIOR OF ROUNDER IS
	COMPONENT REGN_EN_FP IS
		GENERIC ( N : INTEGER:=24);
		PORT (	R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				ENABLE, CLOCK, RESETN : IN STD_LOGIC;
				Q :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;

	SIGNAL ROUND, ZEROS:  STD_LOGIC_VECTOR(N_IN-1 DOWNTO 0);
	SIGNAL IN_REGISTER :STD_LOGIC_VECTOR (M_OUT-1 DOWNTO 0);
BEGIN	
	-- CREAZIONE DEL VETTORE DI ARROTONDAMENTO 'HALF-UP'
	ZEROS (N_IN-1 DOWNTO N_IN-M_OUT)<= (OTHERS=>'0') ;
	ZEROS (N_IN-M_OUT-1)<= '1' ;
	ZEROS (N_IN-M_OUT-2 DOWNTO 0)<= (OTHERS=>'0') ;
	-- ESECUZIONE ARROTONDAMENTO 'TO HALF-UP'
	ROUND <= STD_LOGIC_VECTOR(SIGNED(INPUT) + SIGNED(ZEROS));
	-- USCITA DEL VALORE ARROTONDATO
	IN_REGISTER<= ROUND(N_IN-1 DOWNTO (N_IN-M_OUT));
	REG1: REGN_EN_FP 	GENERIC MAP (M_OUT)
							PORT MAP(IN_REGISTER, '1', CLOCK, RESETN, OUTPUT);
END BEHAVIOR;
