LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TB_BUTTERFLY_singolo IS
END ENTITY;

ARCHITECTURE BEHAVIORAL OF TB_BUTTERFLY_singolo IS
	COMPONENT BUTTERFLY IS
		GENERIC (N: INTEGER:=24);
		PORT (A, B, Wr, Wi  		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				START, CLOCK, RST_n	: IN STD_LOGIC;
				A_O, B_O      		: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0);
				DONE			  		: OUT STD_LOGIC);
	END COMPONENT;
	SIGNAL A, B, Wr, Wi  		: STD_LOGIC_VECTOR(23 DOWNTO 0);
	SIGNAL START, CLOCK, RST_n	: STD_LOGIC;
	SIGNAL A_O, B_O      		: STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL DONE			  		   : STD_LOGIC;
BEGIN
	DUT: BUTTERFLY PORT MAP (A, B, Wr, Wi, START, CLOCK, RST_n, A_O, B_O, DONE);
	
	Wr<="111110100011100111101111"; --0,99999988079071044921875
	Wi<="001110100000011101011111"; --0
	CLK: PROCESS
	BEGIN
		CLOCK<='1';
		WAIT FOR 50 PS;
		CLOCK<='0';
		WAIT FOR 50 PS;
	END PROCESS;
	
	RST: PROCESS
	BEGIN
		RST_n<='0';
		WAIT FOR 130 PS;
		RST_n<='1';
		WAIT;
	END PROCESS;
	
	DATA: PROCESS
	BEGIN
		WAIT FOR 210 PS;
		START<='1';
		WAIT FOR 100 PS;
		START<='0';
		A<="101110001000110001011000"; --  -0.5582
		B<="110001110000001101010011"; --  -0.4452
		WAIT FOR 100 PS;
		A<="110011101001010000101101"; --    -0.3861
		B<="110100010010110000011111"; --     -0.3658
		WAIT;
	END PROCESS;
	-- OUTA=  1372271/2^23 =  0,16358745098114013671875
	-- OUTB= -1372272/2^23 = -0,1635875701904296875
END BEHAVIORAL;