LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX2TO1 IS
GENERIC ( N : INTEGER:=24);
	PORT (I0,I1: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  S	    : IN STD_LOGIC;
		  O     : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY MUX2TO1;

ARCHITECTURE STRUCTURE OF MUX2TO1 IS
BEGIN
O <=	I0 WHEN S='0' ELSE
		I1 WHEN S='1';
END STRUCTURE;