LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SHIFTER IS
	GENERIC ( N: INTEGER:=24;
				 REG_NUM: INTEGER:=2); 
	PORT (	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				EN_SHIFT, CLOCK, RESETN: IN STD_LOGIC;
				OUTPUT :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END SHIFTER;

ARCHITECTURE BEHAVIOR OF SHIFTER IS
	TYPE SHIFT_ARRAY IS ARRAY(0 TO REG_NUM) OF STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	COMPONENT REGN_EN_FP IS
		GENERIC ( N : INTEGER:=24); 
		PORT (	R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				ENABLE, CLOCK, RESETN : IN STD_LOGIC;
				Q :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;
	SIGNAL SHIFT: SHIFT_ARRAY;
BEGIN	
	SHIFT(0)<=STD_LOGIC_VECTOR(A);
	OUTPUT<=(SHIFT(REG_NUM));
	
	GEN_REG: FOR I IN 0 TO REG_NUM-1 GENERATE
      REGX : REGN_EN_FP GENERIC MAP (N)
								PORT MAP(SHIFT(I), EN_SHIFT, CLOCK, RESETN, SHIFT(I+1));
	END GENERATE GEN_REG;
	
END BEHAVIOR;
