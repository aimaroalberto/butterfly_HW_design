LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REGISTER_FILE IS
	GENERIC (N: INTEGER:=24);
	PORT (I0, I1        : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			A_I0, A_I1    : IN STD_LOGIC;--_VECTOR(1 DOWNTO 0);
			WR, CLK, RST_N: IN STD_LOGIC;
			A_O0, A_O1    : IN STD_LOGIC;--_VECTOR(1 DOWNTO 0);
			O0, O1        : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0));
END ENTITY REGISTER_FILE;

ARCHITECTURE BEHAVIORAL OF REGISTER_FILE IS
	TYPE REG_FILE IS ARRAY (0 TO 3) OF STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	SIGNAL I_RF, Q_RF: REG_FILE;
	SIGNAL O_0, O_1: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	SIGNAL EN_R: STD_LOGIC_VECTOR(0 TO 3);
	
	COMPONENT REGN_EN_FP IS
		GENERIC ( N : INTEGER:=24);
		PORT (	R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
					ENABLE, CLOCK, RESETN : IN STD_LOGIC;
					Q :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT REGN_EN_FP;
	
	COMPONENT MUX2TO1 IS
		GENERIC (N : INTEGER:=24);
		PORT 	(	I0,I1: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
					S	  : IN STD_LOGIC;
					O    : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT MUX2TO1;
BEGIN
	O0 <= O_0;
	O1 <= O_1;
	R0: REGN_EN_FP PORT MAP (I_RF(0), EN_R(0), CLK, RST_N, Q_RF(0));
	R1: REGN_EN_FP PORT MAP (I_RF(1), EN_R(1), CLK, RST_N, Q_RF(1));
	R2: REGN_EN_FP PORT MAP (I_RF(2), EN_R(2), CLK, RST_N, Q_RF(2));
	R3: REGN_EN_FP PORT MAP (I_RF(3), EN_R(3), CLK, RST_N, Q_RF(3));
	EN_R(0)<=NOT(A_I0) AND WR;
	EN_R(1)<=(A_I0) AND WR;
	EN_R(2)<=NOT(A_I1) AND WR;
	EN_R(3)<=(A_I1) AND WR;
	I_RF(0)<=I0;
	I_RF(2)<=I1;
	I_RF(1)<=I0;
	I_RF(3)<=I1;
	MUX_0: MUX2TO1 PORT MAP (Q_RF(0), Q_RF(1), A_O0, O_0);
	MUX_1: MUX2TO1 PORT MAP (Q_RF(2), Q_RF(3), A_O1, O_1);

END BEHAVIORAL;