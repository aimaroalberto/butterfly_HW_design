LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ADDER IS
	GENERIC ( N: INTEGER:=24); --dimensione generica
	PORT (	A : IN SIGNED(N-1 DOWNTO 0);
				B : IN SIGNED(N-1 DOWNTO 0);
				EN, CLOCK, RESETN, OP: IN STD_LOGIC;
				OUTPUT :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ADDER;

ARCHITECTURE BEHAVIOR OF ADDER IS
	COMPONENT REGN_EN_FP IS
		GENERIC ( N : INTEGER:=24); --dimensione generica
		PORT (	R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				ENABLE, CLOCK, RESETN : IN STD_LOGIC;
				Q :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;

	SIGNAL E1:  SIGNED(N-1 DOWNTO 0);
	SIGNAL E2,E3:  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	SIGNAL EN_0,EN_1: STD_LOGIC_VECTOR(0 DOWNTO 0);
BEGIN	

	EN_0(0)<=EN;
	-- STADIO DI INGRESSO
	REG1: REGN_EN_FP 	GENERIC MAP (N)
							PORT MAP(STD_LOGIC_VECTOR(E1), EN_0(0), CLOCK, RESETN, E2);
	FF1:  REGN_EN_FP 	GENERIC MAP (1)								
							PORT MAP(EN_0, '1', CLOCK, RESETN, EN_1);
	-- PRIMO LIVELLO DI PIPELINE
	REG2: REGN_EN_FP 	GENERIC MAP (N)
							PORT MAP(E2, EN_1(0), CLOCK, RESETN, E3);
	OUTPUT <= E3;
	E1<= A+B WHEN OP='0' ELSE
		  A-B WHEN OP='1';
END BEHAVIOR;
