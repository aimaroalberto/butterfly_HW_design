LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_3TO1 IS
GENERIC (N:INTEGER:=4);
PORT(	I1: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		I2: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		I3: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		S: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		F: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END MUX_3TO1;

ARCHITECTURE BEHAVIOR OF MUX_3TO1 IS
BEGIN

    F <= I1 WHEN (S = "00") ELSE
         I2 WHEN (S = "01") ELSE
         I3 WHEN (S = "10") ELSE
         "0000";

END BEHAVIOR;