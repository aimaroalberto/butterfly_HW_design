LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MICRO_ROM IS
GENERIC (N : INTEGER := 23; -- NUMBER OF BITS PER ROM WORD
		 M : INTEGER := 4); -- 2^ADDR_BITS = NUMBER OF WORDS IN ROM
PORT (ADDRESS : IN STD_LOGIC_VECTOR(M-1 DOWNTO 0);
	DATA_OUT : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END MICRO_ROM;

ARCHITECTURE BEHAVIORAL OF MICRO_ROM IS
TYPE ROM_TYPE IS ARRAY (2**M-1 DOWNTO 0 ) OF STD_LOGIC_VECTOR (N-1 DOWNTO 0);
SIGNAL ROM : ROM_TYPE;
BEGIN
		ROM(0) <= "10000000000000000000000";
		ROM(1) <= "00111001000000000000000";
		ROM(2) <= "00001010110000000100000";
		ROM(3) <= "00000010000000000100000";
		ROM(4) <= "00000000000000000100010";
		ROM(5) <= "00111101011010000110000";
		ROM(6) <= "00001010111001000110000";
		ROM(7) <= "00000010000000000111000";
		ROM(8) <= "00000000000000000110010";
		ROM(9) <= "00111101011110000110100";
		ROM(10)<= "00001010111001010110100";
		ROM(11)<= "00000010000000110111000";
		ROM(12)<= "00000000000000101110011";
		ROM(13)<= "01111101011110011110100";	
		ROM(14)<= "10000000000000000000000";
		ROM(15)<= "10000000000000000000000";	
					
DATA_OUT <= ROM(CONV_INTEGER(UNSIGNED(ADDRESS)));
END BEHAVIORAL;