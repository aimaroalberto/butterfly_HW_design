LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BUTTERFLY IS
	GENERIC (N: INTEGER:=24);
	PORT (A, B, Wr, Wi  		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			START, CLOCK, RST_n	: IN STD_LOGIC;
			A_O, B_O      		: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0);
			DONE			  		: OUT STD_LOGIC);
END ENTITY BUTTERFLY;

ARCHITECTURE BEHAVIORAL OF BUTTERFLY IS
	COMPONENT CONTROL_UNIT IS
		PORT (	CLOCK,RESET_N : IN STD_LOGIC;
				START, START_R: IN STD_LOGIC;
				INSTRUCTION : OUT STD_LOGIC_VECTOR(20 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT ROUNDER IS
		GENERIC (N_IN : INTEGER := 49;
					M_OUT: INTEGER :=24);
		PORT (	INPUT : IN STD_LOGIC_VECTOR(N_IN-1 DOWNTO 0);
					CLOCK, RESETN : IN STD_LOGIC;
					OUTPUT: OUT STD_LOGIC_VECTOR(M_OUT-1 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT REGN_EN_FP IS
		GENERIC ( N : INTEGER:=24); --dimensione generica
		PORT (	R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
					ENABLE, CLOCK, RESETN : IN STD_LOGIC;
					Q :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT REGN_EN_FP;
	
	COMPONENT MUX2TO1 IS
		GENERIC (N : INTEGER:=24);
		PORT 	(	I0,I1: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
					S	  : IN STD_LOGIC;
					O    : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT MUX2TO1;
	
	COMPONENT SHIFTER IS
		GENERIC ( N: INTEGER:=24;
					 REG_NUM: INTEGER:=2); --dimensione generica
		PORT (	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
					EN_SHIFT, CLOCK, RESETN: IN STD_LOGIC;
					OUTPUT :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT MULTIPLIER IS
		GENERIC ( N, M : INTEGER:=24); --dimensione generica
		PORT (	A : IN SIGNED(N-1 DOWNTO 0);
					B : IN SIGNED(M-1 DOWNTO 0);
					EN, CLOCK, RESETN : IN STD_LOGIC;
					OUTPUT :	OUT STD_LOGIC_VECTOR(M+N-2 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT ADDER IS
		GENERIC ( N: INTEGER:=49); --dimensione generica
		PORT (	A : IN SIGNED(N-1 DOWNTO 0);
					B : IN SIGNED(N-1 DOWNTO 0);
					EN, CLOCK, RESETN, OP: IN STD_LOGIC;
					OUTPUT :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT REGISTER_FILE IS
		GENERIC (N: INTEGER:=24);
		PORT (I0, I1        : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				A_I0, A_I1    : IN STD_LOGIC;--_VECTOR(1 DOWNTO 0);
				WR, CLK, RST_n: IN STD_LOGIC;
				A_O0, A_O1    : IN STD_LOGIC;--_VECTOR(1 DOWNTO 0);
				O0, O1        : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0));
	END COMPONENT;
	
	SIGNAL 	EN_Wr, EN_Wi, Ain, Bin, WR_RF, Aout, Bout, Wout,
				EN_2Ar,EN_2Ai,S2_IN, M, S1_IN, S1, OP1, S2,
				ROUND_B_An, EN_SH_A, EN_B, EN_SH_START: STD_LOGIC;
	SIGNAL	Wr_S, Wi_S, A_S, B_S, W_mul, ROUNDED: STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL	TWO_Ar, TWO_Ai, TWO_A, TWO_A_S: STD_LOGIC_VECTOR(24 DOWNTO 0);
	SIGNAL	O_M: STD_LOGIC_VECTOR(46 DOWNTO 0);
	SIGNAL	O_S1, MUX_S1, S_IN_MUX0, S_IN_MUX1, O_S2, TWO_A_EXT, ROUNDING: STD_LOGIC_VECTOR(48 DOWNTO 0);
	SIGNAL	START_S, START_SH: STD_LOGIC_VECTOR(0 DOWNTO 0);
	SIGNAL	INSTRUCTION : STD_LOGIC_VECTOR(20 DOWNTO 0);
BEGIN
-- -------------------------------------------------------------------------------------------------------------
-- -------------------------------------------------DATAPATH----------------------------------------------------
-- -------------------------------------------------------------------------------------------------------------
	START_S(0)<=START;
	
		REG_WR: REGN_EN_FP 	GENERIC MAP(24)
									PORT MAP (Wr, EN_Wr, CLOCK, RST_n, Wr_S);
		REG_WI: REGN_EN_FP 	GENERIC MAP(24)
									PORT MAP (Wi, EN_Wi, CLOCK, RST_n, Wi_S);
		REG_FILE: REGISTER_FILE 	GENERIC MAP (24)
											PORT MAP (A, B, Ain, Bin, WR_RF, CLOCK, RST_n, Aout, Bout, A_S, B_S);
		MUX_W: MUX2TO1	GENERIC MAP(24)
							PORT MAP(Wi_S, Wr_S, Wout, W_mul);
	-- MOLTIPLICAZIONE PER 2 DI A
	TWO_A_S<= A_S & '0';
	
		REG_2AR: REGN_EN_FP 	GENERIC MAP(25)
									PORT MAP (TWO_A_S, EN_2Ar, CLOCK, RST_n, TWO_Ar);
		REG_2AI: REGN_EN_FP 	GENERIC MAP(25)
									PORT MAP (TWO_A_S, EN_2Ai, CLOCK, RST_n, TWO_Ai);
		MUX_2A: MUX2TO1 	GENERIC MAP (25)
								PORT MAP (TWO_Ai, TWO_Ar, S2_IN, TWO_A);
		MULT: MULTIPLIER  PORT MAP (SIGNED(W_mul),SIGNED(B_S), M, CLOCK, RST_n, O_M);
	-- ALLUNGAMENTO DI SEGNO E RISCALAMENTO DI A
	MUX_S1(48 DOWNTO 23)<= A_S(23)&A_S(23)&  A_S;
	MUX_S1(22 DOWNTO 0) <= (OTHERS=>'0');
	
		S1_MUX: MUX2TO1 	GENERIC MAP (49)
								PORT MAP (O_S1, MUX_S1, S1_IN, S_IN_MUX1);
	-- ALLUNGAMENTO DI SEGNO DELL'USCITA DEL MOLTIPLICATORE						
	S_IN_MUX0<=O_M(46) & O_M(46) & O_M ;
	
		ADD1: ADDER	PORT MAP (SIGNED(S_IN_MUX1), SIGNED(S_IN_MUX0), S1, CLOCK, RST_n, OP1, O_S1);
	-- ALLUNGAMENTO DI SEGNO E RISCALAMENTO DI 2A
	TWO_A_EXT(48 DOWNTO 23)<= TWO_A(24)& TWO_A;
	TWO_A_EXT(22 DOWNTO 0) <= (OTHERS=>'0');
	
		ADD2: ADDER PORT MAP (SIGNED(TWO_A_EXT), SIGNED(O_S1), S2, CLOCK, RST_n, '1', O_S2);
		MUX_ROUND: MUX2TO1	GENERIC MAP(49)
									PORT MAP(O_S1,O_S2,ROUND_B_An, ROUNDING);
		ROUND: ROUNDER	GENERIC MAP(49, 24)
							PORT MAP (ROUNDING, CLOCK, RST_n, ROUNDED);
		SHIFT_A: SHIFTER 	GENERIC MAP (24, 2)
								PORT MAP (ROUNDED, EN_SH_A, CLOCK, RST_n, A_O);
		REG_B_O: REGN_EN_FP 	GENERIC MAP(24)
									PORT MAP (ROUNDED, EN_B, CLOCK, RST_n, B_O);
		SHIFT_START: SHIFTER GENERIC MAP (1, 3)
									PORT MAP(START_S, EN_SH_START, CLOCK, RST_n, START_SH);
		
		CU: CONTROL_UNIT PORT MAP (CLOCK, RST_n, START_S(0), START_SH(0), INSTRUCTION);

-- -------------------------------------------------------------------------------------------------------------
-- --------------------------------ASSOCIAZIONE USCITE A REGISTRO uROM------------------------------------------
-- -------------------------------------------------------------------------------------------------------------
	Ain 		<= INSTRUCTION(20);	
	Bin 		<= INSTRUCTION(19);	
	WR_RF 		<= INSTRUCTION(18);	
	Aout 		<= INSTRUCTION(17);	
	Bout 		<= INSTRUCTION(16);	
	EN_Wr 		<= INSTRUCTION(15);	
	EN_Wi 		<= INSTRUCTION(14);	
	Wout 		<= INSTRUCTION(13);	
	S1_IN 		<= INSTRUCTION(12);	
	S2_IN 		<= INSTRUCTION(11);	
	EN_2Ar 		<= INSTRUCTION(10);	
	EN_2Ai 		<= INSTRUCTION(9);	
	ROUND_B_An 	<= INSTRUCTION(8);	
	EN_SH_A		<= INSTRUCTION(7);
	EN_B 		<= INSTRUCTION(6);	
	M 			<= INSTRUCTION(5);	
	S1 			<= INSTRUCTION(4);	
	OP1			<= INSTRUCTION(3);
	S2 			<= INSTRUCTION(2);
	EN_SH_START	<= INSTRUCTION(1);
	DONE 		<= INSTRUCTION(0);

END BEHAVIORAL;