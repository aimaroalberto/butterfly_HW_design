LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.NUMERIC_STD.ALL;


entity TB_CONTROL_UNIT is

END TB_CONTROL_UNIT;

architecture BEHAVIOR of TB_CONTROL_UNIT is

COMPONENT CONTROL_UNIT is
PORT (	CLOCK,RESET : IN STD_LOGIC;
	    START: IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		INSTRUCTION : OUT STD_LOGIC_VECTOR(22 DOWNTO 0));
END COMPONENT;

	SIGNAL INSTRUCT_OUT: STD_LOGIC_VECTOR(22 DOWNTO 0);
	SIGNAL CLOCK,RESET: STD_LOGIC;
	SIGNAL START: STD_LOGIC_VECTOR (0 DOWNTO 0);
	

BEGIN
DUT: CONTROL_UNIT PORT MAP (CLOCK,RESET,START,INSTRUCT_OUT);
CLK: PROCESS
	BEGIN
		CLOCK<='0';
		WAIT FOR 50 PS;
		CLOCK<='1';
		WAIT FOR 50 PS;
END PROCESS;

ST: PROCESS
	BEGIN
		START<="0";
		WAIT FOR 150 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT FOR 300 PS;
		START<="1";
		WAIT FOR 100 PS;
		START<="0";
		WAIT;
END PROCESS;
	
RST: PROCESS
	BEGIN
		RESET<='0';
		WAIT FOR 25 PS;
		RESET<='1';
		WAIT;
END PROCESS;

END BEHAVIOR;

